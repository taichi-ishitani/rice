module rice_core (
  input var           i_clk,
  input var           i_rst_n,
  rice_bus_if.master  inst_bus_if,
  rice_bus_if.master  data_bus_if
);
endmodule
