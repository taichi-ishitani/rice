typedef tue_status  tb_rice_env_status_base;
