package tb_rice_riscv_pkg;
  import  uvm_pkg::*;

  `include  "uvm_macros.svh"

  typedef enum bit [6:0] {
    TB_RICE_RISCV_OPCODE_BRANCH   = 7'b11_000_11,
    TB_RICE_RISCV_OPCODE_JALR     = 7'b11_001_11,
    TB_RICE_RISCV_OPCODE_JAL      = 7'b11_011_11,
    TB_RICE_RISCV_OPCODE_SYSTEM   = 7'b11_100_11,
    TB_RICE_RISCV_OPCODE_STORE    = 7'b01_000_11,
    TB_RICE_RISCV_OPCODE_OP       = 7'b01_100_11,
    TB_RICE_RISCV_OPCODE_LUI      = 7'b01_101_11,
    TB_RICE_RISCV_OPCODE_LOAD     = 7'b00_000_11,
    TB_RICE_RISCV_OPCODE_MISC_MEM = 7'b00_011_11,
    TB_RICE_RISCV_OPCODE_OP_IMM   = 7'b00_100_11,
    TB_RICE_RISCV_OPCODE_AUIPC    = 7'b00_101_11
  } tb_rice_riscv_opcode;

  typedef enum {
    TB_RICE_RISCV_INST_R_TYPE,
    TB_RICE_RISCV_INST_I_TYPE,
    TB_RICE_RISCV_INST_S_TYPE,
    TB_RICE_RISCV_INST_B_TYPE,
    TB_RICE_RISCV_INST_U_TYPE,
    TB_RICE_RISCV_INST_J_TYPE
  } tb_rice_riscv_inst_type;

  typedef enum {
    TB_RICE_RISCV_INST_NA,
    TB_RICE_RISCV_INST_LUI,
    TB_RICE_RISCV_INST_AUIPC,
    TB_RICE_RISCV_INST_JAL,
    TB_RICE_RISCV_INST_JALR,
    TB_RICE_RISCV_INST_BEQ,
    TB_RICE_RISCV_INST_BNE,
    TB_RICE_RISCV_INST_BLT,
    TB_RICE_RISCV_INST_BGE,
    TB_RICE_RISCV_INST_BLTU,
    TB_RICE_RISCV_INST_BGEU,
    TB_RICE_RISCV_INST_LB,
    TB_RICE_RISCV_INST_LH,
    TB_RICE_RISCV_INST_LW,
    TB_RICE_RISCV_INST_LBU,
    TB_RICE_RISCV_INST_LHU,
    TB_RICE_RISCV_INST_SB,
    TB_RICE_RISCV_INST_SH,
    TB_RICE_RISCV_INST_SW,
    TB_RICE_RISCV_INST_ADDI,
    TB_RICE_RISCV_INST_SLTI,
    TB_RICE_RISCV_INST_SLTIU,
    TB_RICE_RISCV_INST_XORI,
    TB_RICE_RISCV_INST_ORI,
    TB_RICE_RISCV_INST_ANDI,
    TB_RICE_RISCV_INST_SLLI,
    TB_RICE_RISCV_INST_SRLI,
    TB_RICE_RISCV_INST_SRAI,
    TB_RICE_RISCV_INST_ADD,
    TB_RICE_RISCV_INST_SUB,
    TB_RICE_RISCV_INST_SLL,
    TB_RICE_RISCV_INST_SLT,
    TB_RICE_RISCV_INST_SLTU,
    TB_RICE_RISCV_INST_XOR,
    TB_RICE_RISCV_INST_SRL,
    TB_RICE_RISCV_INST_SRA,
    TB_RICE_RISCV_INST_OR,
    TB_RICE_RISCV_INST_AND,
    TB_RICE_RISCV_INST_FENCE,
    TB_RICE_RISCV_INST_FENCE_I,
    TB_RICE_RISCV_INST_ECALL,
    TB_RICE_RISCV_INST_EBREAK,
    TB_RICE_RISCV_INST_CSRRW,
    TB_RICE_RISCV_INST_CSRRS,
    TB_RICE_RISCV_INST_CSRRC,
    TB_RICE_RISCV_INST_CSRRWI,
    TB_RICE_RISCV_INST_CSRRSI,
    TB_RICE_RISCV_INST_CSRRCI,
    TB_RICE_RISCV_INST_MRET
  } tb_rice_riscv_inst;

  `include  "tb_rice_riscv_inst_item.svh"
endpackage
