package tb_rice_core_test_pkg;
  import  uvm_pkg::*;
  import  tue_pkg::*;
  import  tb_rice_bus_pkg::*;
  import  tb_rice_env_base_pkg::*;
  import  tb_rice_core_env_pkg::*;
  import  tb_riscv_test_pkg::*;

  `include  "uvm_macros.svh"
  `include  "tue_macros.svh"

  `include  "tb_rice_core_test_base.svh"
  `include  "tb_rice_core_riscv_test.svh"
endpackage
